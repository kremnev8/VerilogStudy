
module Pacman(clk, shpos, svpos, rgb);
  
  
  
endmodule