
`ifndef MapData_H
`define MapData_H

module MapData(addr_a, addr_b, out_a, out_b);
  
  input [4:0] addr_a;	
  input [4:0] addr_b;	
  
  output [31:0] out_a;
  output [31:0] out_b;
  
  reg [31:0] bitarray[0:31];
  
  assign out_a = bitarray[addr_a];
  assign out_b = bitarray[addr_b];
  
  initial begin/*{w:32,h:32,bpw:32,count:1}*/
    bitarray['h00] = 32'b11111111111111111111111111111111;
    bitarray['h01] = 32'b11111111111111111111111111111111;
    bitarray['h02] = 32'b11110000000000001100000000000011;
    bitarray['h03] = 32'b11110111101111101101111101111011;
    bitarray['h04] = 32'b11110111101111101101111101111011;
    bitarray['h05] = 32'b11110111101111101101111101111011;
    bitarray['h06] = 32'b11110000000000000000000000000011;
    bitarray['h07] = 32'b11110111101101111111101101111011;
    bitarray['h08] = 32'b11110111101101111111101101111011;
    bitarray['h09] = 32'b11110000001100001100001100000011;
    bitarray['h0A] = 32'b11111111101111101101111101111111;
    bitarray['h0B] = 32'b11111111101111101101111101111111;
    bitarray['h0C] = 32'b11111111101100000000001101111111;
    bitarray['h0D] = 32'b11111111101101110011101101111111;
    bitarray['h0E] = 32'b11111111101101110011101101111111;
    bitarray['h0F] = 32'b11110000000001100001100000000011;
    bitarray['h10] = 32'b11111111101101111111101101111111;
    bitarray['h11] = 32'b11111111101101111111101101111111;
    bitarray['h12] = 32'b11111111101100000000001101111111;
    bitarray['h13] = 32'b11111111101101111111101101111111;
    bitarray['h14] = 32'b11111111101101111111101101111111;
    bitarray['h15] = 32'b11110000000000001100000000000011;
    bitarray['h16] = 32'b11110111101111101101111101111011;
    bitarray['h17] = 32'b11110111101111101101111101111011;
    bitarray['h18] = 32'b11110001100000000000000001100011;
    bitarray['h19] = 32'b11111101101101111111101101101111;
    bitarray['h1A] = 32'b11111101101101111111101101101111;
    bitarray['h1B] = 32'b11110000001100000000001100000011;
    bitarray['h1C] = 32'b11111111111111111111111111111111;
    bitarray['h1D] = 32'b11111111111111111111111111111111;
    bitarray['h1E] = 32'b11111111111111111111111111111111;
    bitarray['h1F] = 32'b11111111111111111111111111111111;
  end
  
endmodule

`endif