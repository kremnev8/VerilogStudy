
`define BLACK 3'd0
`define YELLOW 3'd1
`define RED 3'd2
`define WHITE 3'd3
`define BLUE 3'd4
`define PINK 3'd5
`define CYAN 3'd6
`define ORANGE 3'd7

`define FRAME_RATE 10