
`define BLACK 3'd0
`define YELLOW 3'd1
`define RED 3'd2
`define WHITE 3'd3
`define BLUE 3'd4
`define PINK 3'd5
`define CYAN 3'd6
`define ORANGE 3'd7

`define FRAME_RATE 10


`define PACMAN_POS_X 0
`define PACMAN_POS_Y 1
`define PACMAN_ROT   2
`define PACMAN_TIMER 3 
`define PACMAN_WAIT  4 
`define PACMAN_LIFES 5
  
`define WORLD_POS_X  6
`define WORLD_POS_Y  7

`define BLINKY_POS_X 8
`define BLINKY_POS_Y 9
`define BLINKY_ROT   10
`define BLINKY_TIMER 11
`define BLINKY_WAIT  12 
   
`define FRAME_SYNC   22       
`define PELLET_X 23
`define PELLET_Y 24     
`define PELLET_CLEAR 25
`define PELLET_DATA 35      
`define SCORE 26
`define SCORE_DISP 27
   
`define MAP_DATA 32
`define PLAYER_ROT 33