
module BlinkyBitmap(animState, direction, yin, xin, out);
  
  input animState;
  input [1:0] direction;  
  input [3:0] yin;
  input [3:0] xin;
  output out;
  
  reg [31:0] pacman[0:128];
  
  wire [7:0] caseexpr = {1'b0, direction, animState, yin};
  
  assign out = pacman[caseexpr][xin];
  
  initial begin
    /*{w:16,h:16,bpp:2,brev:1, bpw:32,count:8}*/
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b101001010101101000000000;
    pacman['h03] = 32'b11101011010111101011000000;
    pacman['h04] = 32'b111111111010111111111010000;
    pacman['h05] = 32'b111111111010111111111010000;
    pacman['h06] = 32'b101111101010101111101010000;
    pacman['h07] = 32'b10101010101010101010101010100;
    
    pacman['h08] = 32'b10101010101010101010101010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10100010101000001010100010100;
    pacman['h0E] = 32'b10000000101000001010000000100;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b101001010101101000000000;
    pacman['h03] = 32'b11101011010111101011000000;
    pacman['h04] = 32'b111111111010111111111010000;
    pacman['h05] = 32'b111111111010111111111010000;
    pacman['h06] = 32'b101111101010101111101010000;
    pacman['h07] = 32'b10101010101010101010101010100;
    
    pacman['h08] = 32'b10101010101010101010101010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10101010001010101000101010100;
    pacman['h0E] = 32'b101000000010100000001010000;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b101011111010101011111010000;
    pacman['h05] = 32'b101111111110101111111110000;
    pacman['h06] = 32'b101111110100101111110100000;
    pacman['h07] = 32'b10101111110100101111110100100;
    
    pacman['h08] = 32'b10101011111010101011111010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10100010101000001010100010100;
    pacman['h0E] = 32'b10000000101000001010000000100;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b101011111010101011111010000;
    pacman['h05] = 32'b101111111110101111111110000;
    pacman['h06] = 32'b101111110100101111110100000;
    pacman['h07] = 32'b10101111110100101111110100100;
    
    pacman['h08] = 32'b10101011111010101011111010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10101010001010101000101010100;
    pacman['h0E] = 32'b101000000010100000001010000;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b101010101010101010101010000;
    pacman['h05] = 32'b101111101010101111101010000;
    pacman['h06] = 32'b111111111010111111111010000;
    pacman['h07] = 32'b10111111111010111111111010100;
    
    pacman['h08] = 32'b10111101011010111101011010100;
    pacman['h09] = 32'b10101101001010101101001010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10100010101000001010100010100;
    pacman['h0E] = 32'b10000000101000001010000000100;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b101010101010101010101010000;
    pacman['h05] = 32'b101111101010101111101010000;
    pacman['h06] = 32'b111111111010111111111010000;
    pacman['h07] = 32'b10111111111010111111111010100;
    
    pacman['h08] = 32'b10111101011010111101011010100;
    pacman['h09] = 32'b10101101001010101101001010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10101010001010101000101010100;
    pacman['h0E] = 32'b101000000010100000001010000;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b111110101010111110101010000;
    pacman['h05] = 32'b1111111101011111111101010000;
    pacman['h06] = 32'b1010111101011010111101010000;
    pacman['h07] = 32'b11010111101011010111101010100;
    
    pacman['h08] = 32'b10111110101010111110101010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10100010101000001010100010100;
    pacman['h0E] = 32'b10000000101000001010000000100;
    pacman['h0F] = 32'b0;
    
    pacman['h00] = 32'b0;
    pacman['h01] = 32'b1010101000000000000;
    pacman['h02] = 32'b10101010101010100000000;
    pacman['h03] = 32'b1010101010101010101000000;
    pacman['h04] = 32'b111110101010111110101010000;
    pacman['h05] = 32'b1111111101011111111101010000;
    pacman['h06] = 32'b1010111101011010111101010000;
    pacman['h07] = 32'b11010111101011010111101010100;
    
    pacman['h08] = 32'b10111110101010111110101010100;
    pacman['h09] = 32'b10101010101010101010101010100;
    pacman['h0A] = 32'b10101010101010101010101010100;
    pacman['h0B] = 32'b10101010101010101010101010100;
    pacman['h0C] = 32'b10101010101010101010101010100;
    pacman['h0D] = 32'b10101010001010101000101010100;
    pacman['h0E] = 32'b101000000010100000001010000;
    pacman['h0F] = 32'b0;
    
  end
  
endmodule