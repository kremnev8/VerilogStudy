
`define BLACK 3'd0
`define YELLOW 3'd1
`define RED 3'd2
`define WHITE 3'd3
`define BLUE 3'd4
`define PINK 3'd5
`define CYAN 3'd6
`define ORANGE 3'd7

`define FRAME_RATE 10


`define PACMAN_POS_X 0
`define PACMAN_POS_Y 1
`define PACMAN_ROT   2
`define PACMAN_TIMER 3 
`define PACMAN_WAIT  4 
`define PACMAN_LIFES 5
  
`define WORLD_POS_X  6
`define WORLD_POS_Y  7

`define BLINKY_POS_X 8
`define BLINKY_POS_Y 9
`define BLINKY_ROT   10
`define BLINKY_TIMER 11
`define BLINKY_AI  12 
`define BLINKY_AI_TIMER  13
`define BLINKY_WAIT  14 

`define PINKY_POS_X 15
`define PINKY_POS_Y 16
`define PINKY_ROT   17
`define PINKY_TIMER 18
`define PINKY_AI  19
`define PINKY_AI_TIMER  20
`define PINKY_WAIT  21

`define INKY_POS_X 22
`define INKY_POS_Y 23
`define INKY_ROT   24
`define INKY_TIMER 25
`define INKY_AI  26
`define INKY_AI_TIMER  27 
`define INKY_WAIT  28

`define CLYDE_POS_X 29
`define CLYDE_POS_Y 30
`define CLYDE_ROT   31
`define CLYDE_TIMER 32
`define CLYDE_AI  33
`define CLYDE_AI_TIMER  34 
`define CLYDE_WAIT  35

   
`define FRAME_SYNC   36      
`define PELLET_X 37
`define PELLET_Y 38   
`define PELLET_CLEAR 39
`define DISPLAY_FLAGS 40

`define SCORE 41
`define SCORE_DISP 42
  
`define MAP_DATA 48
`define PLAYER_ROT 49
`define FRAME_COUNT 50
`define PELLET_DATA 51



`define A 5'd0
`define B 5'd1
`define C 5'd2
`define D 5'd3
`define E 5'd4
`define F 5'd5
`define G 5'd6
`define H 5'd7
`define I 5'd8
`define J 5'd9
`define K 5'd10
`define L 5'd11
`define M 5'd12
`define N 5'd13
`define O 5'd14
`define P 5'd15
`define Q 5'd16
`define R 5'd17
`define S 5'd18
`define T 5'd19
`define U 5'd20
`define V 5'd21
`define W 5'd22
`define X 5'd23
`define Y 5'd24
`define Z 5'd25

`define EXCLAIM 5'd26
`define SPACE 5'd27