
`ifndef MapData_H
`define MapData_H

module MapData(addr, bits);
  
  input [4:0] addr;	
  output reg [31:0] bits;	// output (5 bits)
  
  always @(*)
    case (addr)
      5'o00: bits = 32'b00000000000000000000000000000000;
      5'o01: bits = 32'b00000000000000000000000000000000;
      5'o02: bits = 32'b00000000000000000000000000000000;
      5'o03: bits = 32'b00000000000000000000000000000000;
      5'o04: bits = 32'b00000000000000000000000000000000;
      5'o05: bits = 32'b00000000000000000000000000000000;
      5'o06: bits = 32'b00000000000000000000000000000000;
      5'o07: bits = 32'b00000000000000000000000000000000;
      5'o10: bits = 32'b00000000000000000000000000000000;
      5'o11: bits = 32'b00000000000000000000000000000000;
      5'o12: bits = 32'b00000000000000000000000000000000;
      5'o13: bits = 32'b00000000000000000000000000000000;
      5'o14: bits = 32'b00000000000000000000000000000000;
      5'o15: bits = 32'b00000000000000000000000000000000;
      5'o16: bits = 32'b00000000000000000000000000000000;
      5'o17: bits = 32'b00000000000000000000000000000000;
      5'o20: bits = 32'b00000000000000000000000000000000;
      5'o21: bits = 32'b00000000000000000000000000000000;
      5'o22: bits = 32'b00000000000000000000000000000000;
      5'o23: bits = 32'b00000000000000000000000000000000;
      5'o24: bits = 32'b00000000000000000000000000000000;
      5'o25: bits = 32'b00000000000000000000000000000000;
      5'o26: bits = 32'b00000000000000000000000000000000;
      5'o27: bits = 32'b00000000000000000000000000000000;
      5'o30: bits = 32'b00000000000000000000000000000000;
      5'o31: bits = 32'b00000000000000000000000000000000;
      5'o32: bits = 32'b00000000000000000000000000000000;
      5'o33: bits = 32'b00000000000000000000000000000000;
      5'o34: bits = 32'b00000000000000000000000000000000;
      5'o35: bits = 32'b00000000000000000000000000000000;
      5'o36: bits = 32'b00000000000000000000000000000000;
      5'o37: bits = 32'b00000000000000000000000000000000;

      default: bits = 0;
    endcase
endmodule

`endif